module mcu_spi(
    input clk,
    
    input spi_clk,
    input spi_ss,
    input [0:0] spi_mosi,
    output [0:0] spi_miso,
    )
